`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////

module sum_nibble(
input [3:0] a, b,
input c0,
output [3:0] s,
output c4,
wire [3:1] c
    );
 sum_comp bit0 (
        .x({a[0]}),
        .y({b[0]}),
        .z(c0),
        .s({s[0]}),
        .c({c[1]}));
 
 sum_comp bit1 (
        .x({a[1]}),
        .y({b[1]}),
        .z({c[1]}),
        .s({s[1]}),
        .c({c[2]})); 
  sum_comp bit2 (
        .x({a[2]}),
        .y({b[2]}),
        .z({c[2]}),
        .s({s[2]}),
        .c({c[3]}));
  sum_comp bit3 (
        .x({a[3]}),
        .y({b[3]}),
        .z({c[3]}),
        .s({s[3]}),
        .c(c4));          
endmodule
